-- Project: adder
-- Testbench: adder_tb
--
-- Simulates the adder entity using functional verification. Input test vectors
-- are read from a file and passed into the design under test. Output test
-- vectors are read from a file and compared to the received outputs from the
-- design under test.
--
-- This testbench writes a log of all events to a file for further analysis.

library ieee;
use ieee.std_logic_1164.all;

library std;
use std.textio.all;

library veriti;
use veriti.test.all;

library amp;
use amp.prelude.all;

entity adder_tb is
  generic(
    WORD_SIZE: psize := 16
  );
end entity;


architecture sim of adder_tb is
  -- This record is auto-generated by veriti; DO NOT EDIT.
  type adder_bfm is record
    cin: logic;
    in0: logics(WORD_SIZE-1 downto 0);
    in1: logics(WORD_SIZE-1 downto 0);
    sum: logics(WORD_SIZE-1 downto 0);
    cout: logic;
  end record;
    
  signal bfm: adder_bfm;

  signal clk: logic := '0';
  signal halt: bool := false;

  -- Declare internal required testbench signals
  constant TIMEOUT_LIMIT: usize := 1_000;

  file events: text open write_mode is "events.log";
begin
  -- Instantiate the design under test
  dut: entity work.adder
    generic map (
      WORD_SIZE => WORD_SIZE
    ) port map (
      cin  => bfm.cin,
      in0  => bfm.in0,
      in1  => bfm.in1,
      sum  => bfm.sum,
      cout => bfm.cout
    );

  -- Generate a clock for the testbench
  spin_clock(clk, 40 ns, halt);

  -- Test reading a file filled with test vectors
  driver: process
    file inputs: text open read_mode is "inputs.txt";

    -- This procedure is auto-generated by veriti; DO NOT EDIT.
    procedure send_transaction(file fd: text) is
      variable row: line;
    begin
      if endfile(fd) = false then
        readline(fd, row);
        drive(row, bfm.cin);
        drive(row, bfm.in0);
        drive(row, bfm.in1);
      end if;
    end procedure;

  begin  
    -- Drive transactions
    while endfile(inputs) = false loop
      send_transaction(inputs);
      wait until rising_edge(clk);
    end loop;
    -- Wait for all outputs to be checked
    wait;
  end process;

  checker: process
    file outputs: text open read_mode is "outputs.txt";

    -- This procedure is auto-generated by veriti; DO NOT EDIT.
    procedure score_transaction(file fd: text) is 
      variable row: line;
      variable expct: adder_bfm;
    begin
      if endfile(fd) = false then
        readline(fd, row);
        load(row, expct.sum);
        assert_eq(events, bfm.sum, expct.sum, "sum");
        load(row, expct.cout);
        assert_eq(events, bfm.cout, expct.cout, "cout");
      end if;
    end procedure;

  begin
    while endfile(outputs) = false loop
      -- Wait for a valid time to check
      wait until rising_edge(clk);
      -- Compare outputs
      score_transaction(outputs);
    end loop;
    -- Halt the simulation
    complete(halt);
  end process;

end architecture;